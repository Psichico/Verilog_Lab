
module Question4_testbench();

	reg [15:0] in;
	wire [3:0] out;

	Question4 tb1(.in(in),.out(out));
	
	initial begin
	
		in = 16'b0000_0000_0000_0001;
		#10;
		in = 16'b0000_0000_0000_0010;
		#10;
		in = 16'b0000_0000_0000_0100;
		#10;
		in = 16'b0000_0000_0000_1000;
		#10;
		in = 16'b0000_0000_0001_0000;
		#10;
		in = 16'b0000_0000_0010_0000;
		#10;
		in = 16'b0000_0000_0100_0000;
		#10;
		in = 16'b0000_0000_1000_0000;
		#10;
		in = 16'b0000_0001_0000_0000;
		#10;
		in = 16'b0000_0010_0000_0000;
		#10;
		in = 16'b0000_0100_0000_0000;
		#10;
		in = 16'b0000_1000_0000_0000;
		#10;
		in = 16'b0001_0000_0000_0000;
		#10;
		in = 16'b0010_0000_0000_0000;
		#10;
		in = 16'b0100_0000_0000_0000;
		#10;
		in = 16'b1000_0000_0000_0000;
		#10;
		#100;
	
	end

endmodule
